----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    12:45:46 08/02/2015 
-- Design Name: 
-- Module Name:    IntCtrl - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity INTctrl is
    port(
        intr: in std_logic_vector(7 downto 0);
        newImr: in std_logic_vector(7 downto 0);
        intrUpdate: in std_logic;
        imrUpdate: in std_logic;
        isrUpdate: in std_logic;
        entered : in std_logic;
        nextService: out std_logic; -- ����CPU���Խ���
        intServicePort: out integer;
        nowimr: out std_logic_vector(7 downto 0)
    );
end INTctrl;

architecture Behavioral of INTctrl is
	-- signal irr: std_logic_vector(7 downto 0):= "00000000"; -- ����Ӧ�����
	signal isr: std_logic_vector(7 downto 0):= "00000000"; -- ��������ִ�е��жϷ������
	signal imr: std_logic_vector(7 downto 0):= "10000000"; -- ������
    type stackType is array(0 to 8) of integer;
    signal PortStack : stackType := (8, 0, 0, 0, 0, 0, 0, 0, 0);
    signal stackTop : integer := 0;
    signal pushStack, popStack : std_logic := '0';
    signal runningPort : integer := 8;
begin
	intServicePort <= runningPort;
    nowimr <= imr;
    imr <= newImr when rising_edge(imrUpdate);
	
    process(intrUpdate, entered, isrUpdate, intr, isr, imr)
    begin
        if intrUpdate = '1' then
            if intr(0) = '1' and imr(0) = '0' then
                nextService <= '1';
                runningPort <= 0;
            elsif intr(1) = '1' and imr(1) = '0' then
                nextService <= '1';
                runningPort <= 1;
            elsif intr(2) = '1' and imr(2) = '0' then
                nextService <= '1';
                runningPort <= 2;
            elsif intr(3) = '1' and imr(3) = '0' then
                nextService <= '1';
                runningPort <= 3;
            elsif intr(4) = '1' and imr(4) = '0' then
                nextService <= '1';
                runningPort <= 4;
            elsif intr(5) = '1' and imr(5) = '0' then
                nextService <= '1';
                runningPort <= 5;
            elsif intr(6) = '1' and imr(6) = '0' then
                nextService <= '1';
                runningPort <= 6;
            elsif intr(7) = '1' and imr(7) = '0' then
                nextService <= '1';
                runningPort <= 7;
            else
                nextService <= '0';
                runningPort <= 8;
            end if;
        elsif entered = '1' then
            nextService <= '0';
            isr(runningPort) <= '1';
        elsif isrUpdate = '1' and isrUpdate'event then
            isr(runningPort) <= '0';
            runningPort <= 8;
        end if;
    end process;

end Behavioral;